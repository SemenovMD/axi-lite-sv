package axil_pkg;

    // AXI-Lite Master
    parameter   AXI_DATA_WIDTH  = 32;
    parameter   AXI_ADDR_WIDTH  = 32;

endpackage