package axil_pkg;

    parameter                               AXI_DATA_WIDTH                  = 32;
    parameter                               AXI_ADDR_WIDTH                  = 32;

    parameter                               MEMORY_RAM                      = 1024;

endpackage