package axil_pkg;

    parameter                               AXI_DATA_WIDTH                  = 32;
    parameter                               AXI_ADDR_WIDTH                  = 32;

    parameter                               GPIO_DATA_WIDTH                 = 4;

endpackage